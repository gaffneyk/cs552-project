/*
   CS/ECE 552, Spring '19
   Homework #6, Problem #1
  
   This module determines all of the control logic for the processor.
*/
module control (/*AUTOARG*/
                // Outputs
                err, 
                RegDst,
                SESel,
                RegWrite,
                DMemWrite,
                DMemEn,
                ALUSrc2,
                PCSrc,
                PCImm,
                MemToReg,
                DMemDump,
                Jump,
                // Inputs
                OpCode,
                Funct
                );

   // inputs
   input [4:0]  OpCode;
   input [1:0]  Funct;
   
   // outputs
   output       err;
   output       RegWrite, DMemWrite, DMemEn, ALUSrc2, PCSrc, 
                PCImm, MemToReg, DMemDump, Jump;
   output [1:0] RegDst;
   output [2:0] SESel;

   /* YOUR CODE HERE */

errMod errMod1 (.OpCode(OpCode), .Funct(Funct), .err(err));

RegDstMod RegDstMod1 (.OpCode(OpCode), .RegDst(RegDst));
SESelMod SESelMod1 (.OpCode(OpCode), .SESel(SESel));
RegWriteMod RegWriteMod1 (.OpCode(OpCode), .RegWrite(RegWrite));
DMemWriteMod DMemWriteMod1 (.OpCode(OpCode), .DMemWrite(DMemWrite));
DMemEnMod DMemEnMod1 (.OpCode(OpCode), .DMemEn(DMemEn));
ALUSrc2Mod ALUSrc2Mod1 (.OpCode(OpCode), .ALUSrc2(ALUSrc2));
PCSrcMod PCSrcMod1 (.OpCode(OpCode), .PCSrc(PCSrc));
PCImmMod PCImmMod1 (.OpCode(OpCode), .PCImm(PCImm));
MemToRegMod MemToRegMod1 (.OpCode(OpCode), .MemToReg(MemToReg));
DMemDumpMod DMemDumpMod1 (.OpCode(OpCode), .DMemDump(DMemDump));
JumpMod JumpMod1 (.OpCode(OpCode), .Jump(Jump));


endmodule
